package UVInterp;

    import Semi_FIFOF :: *;
    import FIFOF :: *;
    import Reciprocal :: *;
    import Vector :: *;

    typedef struct {
        Vector #(3, Int #(27)) edge_vec;
        Vector #(3, Vector #(2, Int #(27))) uv;
    } UVInterpIn
    deriving (Bits, FShow);

    typedef struct {
        Int #(27) u;
        Int #(27) v;
    } UVInterpOut
    deriving (Bits, FShow);

    interface UVInterp;
        interface FIFOF_I #(UVInterpIn) in;
        interface FIFOF_O #(UVInterpOut) out;
    endinterface

    (* synthesize *)
    module mkUVInterp(UVInterp);
        FIFOF #(UVInterpIn) f_in <- mkFIFOF;
        FIFOF #(UVInterpOut) f_out <- mkFIFOF;

        Reciprocal #(27) reciprocal <- mkReciprocal;
        FIFOF #(Tuple2 #(Vector #(3, Int #(27)), Vector #(3, Int #(27)))) s0 <- mkFIFOF;
        FIFOF #(Tuple2 #(Int #(27), Int #(27))) s1 <- mkFIFOF;

        rule rl_s0;
            let d = f_in.first; f_in.deq;
            let s = d.edge_vec[0] + d.edge_vec[1] + d.edge_vec[2];
            reciprocal.in.enq(pack(s));
            Vector #(3, Int #(27)) u = newVector;
            Vector #(3, Int #(27)) v = newVector;
            for(Integer i = 0; i < 3; i = i + 1) begin
                Int #(54) uu = extend(d.edge_vec[i]) * extend(d.uv[i][0]);
                u[i] = truncate(uu >> 27);
                Int #(54) vv = extend(d.edge_vec[i]) * extend(d.uv[i][1]);
                v[i] = truncate(vv >> 27);
            end
            s0.enq(tuple2(u, v));
        endrule

        rule rl_s1;
            match {.u, .v} = s0.first; s0.deq;
            let uu = u[0] + u[1] + u[2];
            let vv = v[0] + v[1] + v[2];
            s1.enq(tuple2(uu, vv));
        endrule

        rule rl_s2;
            match {.u, .v} = s1.first; s1.deq;
            let w <- pop_o(reciprocal.out);
            Int #(54) u0 = extend(u) * unpack(zeroExtend(w.value));
            Int #(54) v0 = extend(v) * unpack(zeroExtend(w.value));
            Int #(27) u1 = truncate(u0 >> 26 - w.shift);
            Int #(27) v1 = truncate(v0 >> 26 - w.shift);
            f_out.enq(UVInterpOut {u: u1, v: v1});
        endrule

        interface in = to_FIFOF_I(f_in);
        interface out = to_FIFOF_O(f_out);
    endmodule

endpackage